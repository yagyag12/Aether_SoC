VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO aether_soc
  CLASS BLOCK ;
  FOREIGN aether_soc ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 310.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 998.245 406.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 310.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 998.245 560.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 310.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 998.245 713.840 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 310.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 998.245 867.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 202.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 347.485 1174.640 498.715 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 619.640 1174.640 800.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 925.080 1174.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1188.880 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 310.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 998.245 329.840 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 310.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 998.245 483.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 310.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 998.245 637.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 310.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 998.245 790.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 202.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 347.485 1097.840 802.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 923.005 1097.840 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1049.380 187.440 1050.980 362.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1049.380 486.640 1050.980 634.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1049.380 785.840 1050.980 938.640 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 374.990 1196.000 375.270 1200.000 ;
    END
  END clk
  PIN dmem_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END dmem_addr[0]
  PIN dmem_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END dmem_addr[10]
  PIN dmem_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END dmem_addr[11]
  PIN dmem_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END dmem_addr[12]
  PIN dmem_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END dmem_addr[13]
  PIN dmem_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END dmem_addr[14]
  PIN dmem_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END dmem_addr[15]
  PIN dmem_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END dmem_addr[16]
  PIN dmem_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END dmem_addr[17]
  PIN dmem_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END dmem_addr[18]
  PIN dmem_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END dmem_addr[19]
  PIN dmem_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END dmem_addr[1]
  PIN dmem_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END dmem_addr[20]
  PIN dmem_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END dmem_addr[21]
  PIN dmem_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END dmem_addr[22]
  PIN dmem_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END dmem_addr[23]
  PIN dmem_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END dmem_addr[24]
  PIN dmem_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END dmem_addr[25]
  PIN dmem_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END dmem_addr[26]
  PIN dmem_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END dmem_addr[27]
  PIN dmem_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END dmem_addr[28]
  PIN dmem_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END dmem_addr[29]
  PIN dmem_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END dmem_addr[2]
  PIN dmem_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END dmem_addr[30]
  PIN dmem_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END dmem_addr[31]
  PIN dmem_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END dmem_addr[3]
  PIN dmem_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END dmem_addr[4]
  PIN dmem_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END dmem_addr[5]
  PIN dmem_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END dmem_addr[6]
  PIN dmem_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END dmem_addr[7]
  PIN dmem_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END dmem_addr[8]
  PIN dmem_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END dmem_addr[9]
  PIN dmem_ren
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END dmem_ren
  PIN dmem_wdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END dmem_wdata[0]
  PIN dmem_wdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END dmem_wdata[10]
  PIN dmem_wdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END dmem_wdata[11]
  PIN dmem_wdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END dmem_wdata[12]
  PIN dmem_wdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END dmem_wdata[13]
  PIN dmem_wdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END dmem_wdata[14]
  PIN dmem_wdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END dmem_wdata[15]
  PIN dmem_wdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END dmem_wdata[16]
  PIN dmem_wdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END dmem_wdata[17]
  PIN dmem_wdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END dmem_wdata[18]
  PIN dmem_wdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END dmem_wdata[19]
  PIN dmem_wdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END dmem_wdata[1]
  PIN dmem_wdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END dmem_wdata[20]
  PIN dmem_wdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END dmem_wdata[21]
  PIN dmem_wdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END dmem_wdata[22]
  PIN dmem_wdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END dmem_wdata[23]
  PIN dmem_wdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END dmem_wdata[24]
  PIN dmem_wdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END dmem_wdata[25]
  PIN dmem_wdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END dmem_wdata[26]
  PIN dmem_wdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END dmem_wdata[27]
  PIN dmem_wdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END dmem_wdata[28]
  PIN dmem_wdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END dmem_wdata[29]
  PIN dmem_wdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END dmem_wdata[2]
  PIN dmem_wdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END dmem_wdata[30]
  PIN dmem_wdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END dmem_wdata[31]
  PIN dmem_wdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END dmem_wdata[3]
  PIN dmem_wdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END dmem_wdata[4]
  PIN dmem_wdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END dmem_wdata[5]
  PIN dmem_wdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END dmem_wdata[6]
  PIN dmem_wdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END dmem_wdata[7]
  PIN dmem_wdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END dmem_wdata[8]
  PIN dmem_wdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END dmem_wdata[9]
  PIN dmem_wen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END dmem_wen
  PIN dmem_wmask[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END dmem_wmask[0]
  PIN dmem_wmask[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END dmem_wmask[1]
  PIN dmem_wmask[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END dmem_wmask[2]
  PIN dmem_wmask[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END dmem_wmask[3]
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 516.840 1500.000 517.440 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 788.840 1500.000 789.440 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 816.040 1500.000 816.640 ;
    END
  END gpio_in[11]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 544.040 1500.000 544.640 ;
    END
  END gpio_in[1]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 571.240 1500.000 571.840 ;
    END
  END gpio_in[2]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 598.440 1500.000 599.040 ;
    END
  END gpio_in[3]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 625.640 1500.000 626.240 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 652.840 1500.000 653.440 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 680.040 1500.000 680.640 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 707.240 1500.000 707.840 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 734.440 1500.000 735.040 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 761.640 1500.000 762.240 ;
    END
  END gpio_in[9]
  PIN gpio_led[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 408.040 1500.000 408.640 ;
    END
  END gpio_led[0]
  PIN gpio_led[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 435.240 1500.000 435.840 ;
    END
  END gpio_led[1]
  PIN gpio_led[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 462.440 1500.000 463.040 ;
    END
  END gpio_led[2]
  PIN gpio_led[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 489.640 1500.000 490.240 ;
    END
  END gpio_led[3]
  PIN gpio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 843.240 1500.000 843.840 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1115.240 1500.000 1115.840 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1142.440 1500.000 1143.040 ;
    END
  END gpio_out[11]
  PIN gpio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 870.440 1500.000 871.040 ;
    END
  END gpio_out[1]
  PIN gpio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 897.640 1500.000 898.240 ;
    END
  END gpio_out[2]
  PIN gpio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 924.840 1500.000 925.440 ;
    END
  END gpio_out[3]
  PIN gpio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 952.040 1500.000 952.640 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 979.240 1500.000 979.840 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1006.440 1500.000 1007.040 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1033.640 1500.000 1034.240 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1060.840 1500.000 1061.440 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1088.040 1500.000 1088.640 ;
    END
  END gpio_out[9]
  PIN gpio_sw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 299.240 1500.000 299.840 ;
    END
  END gpio_sw[0]
  PIN gpio_sw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 326.440 1500.000 327.040 ;
    END
  END gpio_sw[1]
  PIN gpio_sw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 353.640 1500.000 354.240 ;
    END
  END gpio_sw[2]
  PIN gpio_sw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 380.840 1500.000 381.440 ;
    END
  END gpio_sw[3]
  PIN imem_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END imem_addr[0]
  PIN imem_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END imem_addr[10]
  PIN imem_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END imem_addr[11]
  PIN imem_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END imem_addr[12]
  PIN imem_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END imem_addr[13]
  PIN imem_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END imem_addr[14]
  PIN imem_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END imem_addr[15]
  PIN imem_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END imem_addr[16]
  PIN imem_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END imem_addr[17]
  PIN imem_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END imem_addr[18]
  PIN imem_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END imem_addr[19]
  PIN imem_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END imem_addr[1]
  PIN imem_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END imem_addr[20]
  PIN imem_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END imem_addr[21]
  PIN imem_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END imem_addr[22]
  PIN imem_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END imem_addr[23]
  PIN imem_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END imem_addr[24]
  PIN imem_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END imem_addr[25]
  PIN imem_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END imem_addr[26]
  PIN imem_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END imem_addr[27]
  PIN imem_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END imem_addr[28]
  PIN imem_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END imem_addr[29]
  PIN imem_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END imem_addr[2]
  PIN imem_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END imem_addr[30]
  PIN imem_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END imem_addr[31]
  PIN imem_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END imem_addr[3]
  PIN imem_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END imem_addr[4]
  PIN imem_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END imem_addr[5]
  PIN imem_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END imem_addr[6]
  PIN imem_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END imem_addr[7]
  PIN imem_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END imem_addr[8]
  PIN imem_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END imem_addr[9]
  PIN imem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END imem_rdata[0]
  PIN imem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END imem_rdata[10]
  PIN imem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END imem_rdata[11]
  PIN imem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END imem_rdata[12]
  PIN imem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END imem_rdata[13]
  PIN imem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END imem_rdata[14]
  PIN imem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END imem_rdata[15]
  PIN imem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END imem_rdata[16]
  PIN imem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END imem_rdata[17]
  PIN imem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END imem_rdata[18]
  PIN imem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END imem_rdata[19]
  PIN imem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END imem_rdata[1]
  PIN imem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END imem_rdata[20]
  PIN imem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END imem_rdata[21]
  PIN imem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END imem_rdata[22]
  PIN imem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END imem_rdata[23]
  PIN imem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.561499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END imem_rdata[24]
  PIN imem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END imem_rdata[25]
  PIN imem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END imem_rdata[26]
  PIN imem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 8.259300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END imem_rdata[27]
  PIN imem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.128699 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END imem_rdata[28]
  PIN imem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END imem_rdata[29]
  PIN imem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.563399 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END imem_rdata[2]
  PIN imem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END imem_rdata[30]
  PIN imem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END imem_rdata[31]
  PIN imem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.563399 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END imem_rdata[3]
  PIN imem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.171599 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END imem_rdata[4]
  PIN imem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.955200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END imem_rdata[5]
  PIN imem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 8.694000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END imem_rdata[6]
  PIN imem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END imem_rdata[7]
  PIN imem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END imem_rdata[8]
  PIN imem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END imem_rdata[9]
  PIN pwm_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1169.640 1500.000 1170.240 ;
    END
  END pwm_out
  PIN ram_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END ram_rdata[0]
  PIN ram_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END ram_rdata[10]
  PIN ram_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END ram_rdata[11]
  PIN ram_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END ram_rdata[12]
  PIN ram_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END ram_rdata[13]
  PIN ram_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END ram_rdata[14]
  PIN ram_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END ram_rdata[15]
  PIN ram_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END ram_rdata[16]
  PIN ram_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END ram_rdata[17]
  PIN ram_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END ram_rdata[18]
  PIN ram_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END ram_rdata[19]
  PIN ram_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END ram_rdata[1]
  PIN ram_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END ram_rdata[20]
  PIN ram_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END ram_rdata[21]
  PIN ram_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END ram_rdata[22]
  PIN ram_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END ram_rdata[23]
  PIN ram_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END ram_rdata[24]
  PIN ram_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END ram_rdata[25]
  PIN ram_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END ram_rdata[26]
  PIN ram_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END ram_rdata[27]
  PIN ram_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END ram_rdata[28]
  PIN ram_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END ram_rdata[29]
  PIN ram_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END ram_rdata[2]
  PIN ram_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END ram_rdata[30]
  PIN ram_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END ram_rdata[31]
  PIN ram_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END ram_rdata[3]
  PIN ram_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END ram_rdata[4]
  PIN ram_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END ram_rdata[5]
  PIN ram_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END ram_rdata[6]
  PIN ram_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END ram_rdata[7]
  PIN ram_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END ram_rdata[8]
  PIN ram_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END ram_rdata[9]
  PIN ram_rvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END ram_rvalid
  PIN rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 1124.790 1196.000 1125.070 1200.000 ;
    END
  END rstn
  PIN spi_clk
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 81.640 1500.000 82.240 ;
    END
  END spi_clk
  PIN spi_master_cs[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 190.440 1500.000 191.040 ;
    END
  END spi_master_cs[0]
  PIN spi_master_cs[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 217.640 1500.000 218.240 ;
    END
  END spi_master_cs[1]
  PIN spi_master_cs[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 244.840 1500.000 245.440 ;
    END
  END spi_master_cs[2]
  PIN spi_master_cs[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 272.040 1500.000 272.640 ;
    END
  END spi_master_cs[3]
  PIN spi_miso
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 108.840 1500.000 109.440 ;
    END
  END spi_miso
  PIN spi_mosi
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 136.040 1500.000 136.640 ;
    END
  END spi_mosi
  PIN spi_slave_csn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 163.240 1500.000 163.840 ;
    END
  END spi_slave_csn
  PIN uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 27.240 1500.000 27.840 ;
    END
  END uart_rx
  PIN uart_tx
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 54.440 1500.000 55.040 ;
    END
  END uart_tx
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 1494.270 1188.830 ;
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1188.725 ;
      LAYER met1 ;
        RECT 4.210 10.640 1494.080 1188.880 ;
      LAYER met2 ;
        RECT 4.230 1195.720 374.710 1196.530 ;
        RECT 375.550 1195.720 1124.510 1196.530 ;
        RECT 1125.350 1195.720 1492.610 1196.530 ;
        RECT 4.230 10.695 1492.610 1195.720 ;
      LAYER met3 ;
        RECT 3.990 1170.640 1496.000 1188.805 ;
        RECT 3.990 1169.240 1495.600 1170.640 ;
        RECT 3.990 1163.840 1496.000 1169.240 ;
        RECT 4.400 1162.440 1496.000 1163.840 ;
        RECT 3.990 1157.040 1496.000 1162.440 ;
        RECT 4.400 1155.640 1496.000 1157.040 ;
        RECT 3.990 1150.240 1496.000 1155.640 ;
        RECT 4.400 1148.840 1496.000 1150.240 ;
        RECT 3.990 1143.440 1496.000 1148.840 ;
        RECT 4.400 1142.040 1495.600 1143.440 ;
        RECT 3.990 1136.640 1496.000 1142.040 ;
        RECT 4.400 1135.240 1496.000 1136.640 ;
        RECT 3.990 1129.840 1496.000 1135.240 ;
        RECT 4.400 1128.440 1496.000 1129.840 ;
        RECT 3.990 1123.040 1496.000 1128.440 ;
        RECT 4.400 1121.640 1496.000 1123.040 ;
        RECT 3.990 1116.240 1496.000 1121.640 ;
        RECT 4.400 1114.840 1495.600 1116.240 ;
        RECT 3.990 1109.440 1496.000 1114.840 ;
        RECT 4.400 1108.040 1496.000 1109.440 ;
        RECT 3.990 1102.640 1496.000 1108.040 ;
        RECT 4.400 1101.240 1496.000 1102.640 ;
        RECT 3.990 1095.840 1496.000 1101.240 ;
        RECT 4.400 1094.440 1496.000 1095.840 ;
        RECT 3.990 1089.040 1496.000 1094.440 ;
        RECT 4.400 1087.640 1495.600 1089.040 ;
        RECT 3.990 1082.240 1496.000 1087.640 ;
        RECT 4.400 1080.840 1496.000 1082.240 ;
        RECT 3.990 1075.440 1496.000 1080.840 ;
        RECT 4.400 1074.040 1496.000 1075.440 ;
        RECT 3.990 1068.640 1496.000 1074.040 ;
        RECT 4.400 1067.240 1496.000 1068.640 ;
        RECT 3.990 1061.840 1496.000 1067.240 ;
        RECT 4.400 1060.440 1495.600 1061.840 ;
        RECT 3.990 1055.040 1496.000 1060.440 ;
        RECT 4.400 1053.640 1496.000 1055.040 ;
        RECT 3.990 1048.240 1496.000 1053.640 ;
        RECT 4.400 1046.840 1496.000 1048.240 ;
        RECT 3.990 1041.440 1496.000 1046.840 ;
        RECT 4.400 1040.040 1496.000 1041.440 ;
        RECT 3.990 1034.640 1496.000 1040.040 ;
        RECT 4.400 1033.240 1495.600 1034.640 ;
        RECT 3.990 1027.840 1496.000 1033.240 ;
        RECT 4.400 1026.440 1496.000 1027.840 ;
        RECT 3.990 1021.040 1496.000 1026.440 ;
        RECT 4.400 1019.640 1496.000 1021.040 ;
        RECT 3.990 1014.240 1496.000 1019.640 ;
        RECT 4.400 1012.840 1496.000 1014.240 ;
        RECT 3.990 1007.440 1496.000 1012.840 ;
        RECT 4.400 1006.040 1495.600 1007.440 ;
        RECT 3.990 1000.640 1496.000 1006.040 ;
        RECT 4.400 999.240 1496.000 1000.640 ;
        RECT 3.990 993.840 1496.000 999.240 ;
        RECT 4.400 992.440 1496.000 993.840 ;
        RECT 3.990 987.040 1496.000 992.440 ;
        RECT 4.400 985.640 1496.000 987.040 ;
        RECT 3.990 980.240 1496.000 985.640 ;
        RECT 4.400 978.840 1495.600 980.240 ;
        RECT 3.990 973.440 1496.000 978.840 ;
        RECT 4.400 972.040 1496.000 973.440 ;
        RECT 3.990 966.640 1496.000 972.040 ;
        RECT 4.400 965.240 1496.000 966.640 ;
        RECT 3.990 959.840 1496.000 965.240 ;
        RECT 4.400 958.440 1496.000 959.840 ;
        RECT 3.990 953.040 1496.000 958.440 ;
        RECT 4.400 951.640 1495.600 953.040 ;
        RECT 3.990 946.240 1496.000 951.640 ;
        RECT 4.400 944.840 1496.000 946.240 ;
        RECT 3.990 939.440 1496.000 944.840 ;
        RECT 4.400 938.040 1496.000 939.440 ;
        RECT 3.990 932.640 1496.000 938.040 ;
        RECT 4.400 931.240 1496.000 932.640 ;
        RECT 3.990 925.840 1496.000 931.240 ;
        RECT 4.400 924.440 1495.600 925.840 ;
        RECT 3.990 919.040 1496.000 924.440 ;
        RECT 4.400 917.640 1496.000 919.040 ;
        RECT 3.990 912.240 1496.000 917.640 ;
        RECT 4.400 910.840 1496.000 912.240 ;
        RECT 3.990 905.440 1496.000 910.840 ;
        RECT 4.400 904.040 1496.000 905.440 ;
        RECT 3.990 898.640 1496.000 904.040 ;
        RECT 4.400 897.240 1495.600 898.640 ;
        RECT 3.990 891.840 1496.000 897.240 ;
        RECT 4.400 890.440 1496.000 891.840 ;
        RECT 3.990 885.040 1496.000 890.440 ;
        RECT 4.400 883.640 1496.000 885.040 ;
        RECT 3.990 878.240 1496.000 883.640 ;
        RECT 4.400 876.840 1496.000 878.240 ;
        RECT 3.990 871.440 1496.000 876.840 ;
        RECT 4.400 870.040 1495.600 871.440 ;
        RECT 3.990 864.640 1496.000 870.040 ;
        RECT 4.400 863.240 1496.000 864.640 ;
        RECT 3.990 857.840 1496.000 863.240 ;
        RECT 4.400 856.440 1496.000 857.840 ;
        RECT 3.990 851.040 1496.000 856.440 ;
        RECT 4.400 849.640 1496.000 851.040 ;
        RECT 3.990 844.240 1496.000 849.640 ;
        RECT 4.400 842.840 1495.600 844.240 ;
        RECT 3.990 837.440 1496.000 842.840 ;
        RECT 4.400 836.040 1496.000 837.440 ;
        RECT 3.990 830.640 1496.000 836.040 ;
        RECT 4.400 829.240 1496.000 830.640 ;
        RECT 3.990 823.840 1496.000 829.240 ;
        RECT 4.400 822.440 1496.000 823.840 ;
        RECT 3.990 817.040 1496.000 822.440 ;
        RECT 4.400 815.640 1495.600 817.040 ;
        RECT 3.990 810.240 1496.000 815.640 ;
        RECT 4.400 808.840 1496.000 810.240 ;
        RECT 3.990 803.440 1496.000 808.840 ;
        RECT 4.400 802.040 1496.000 803.440 ;
        RECT 3.990 796.640 1496.000 802.040 ;
        RECT 4.400 795.240 1496.000 796.640 ;
        RECT 3.990 789.840 1496.000 795.240 ;
        RECT 4.400 788.440 1495.600 789.840 ;
        RECT 3.990 783.040 1496.000 788.440 ;
        RECT 4.400 781.640 1496.000 783.040 ;
        RECT 3.990 776.240 1496.000 781.640 ;
        RECT 4.400 774.840 1496.000 776.240 ;
        RECT 3.990 769.440 1496.000 774.840 ;
        RECT 4.400 768.040 1496.000 769.440 ;
        RECT 3.990 762.640 1496.000 768.040 ;
        RECT 4.400 761.240 1495.600 762.640 ;
        RECT 3.990 755.840 1496.000 761.240 ;
        RECT 4.400 754.440 1496.000 755.840 ;
        RECT 3.990 749.040 1496.000 754.440 ;
        RECT 4.400 747.640 1496.000 749.040 ;
        RECT 3.990 742.240 1496.000 747.640 ;
        RECT 4.400 740.840 1496.000 742.240 ;
        RECT 3.990 735.440 1496.000 740.840 ;
        RECT 4.400 734.040 1495.600 735.440 ;
        RECT 3.990 728.640 1496.000 734.040 ;
        RECT 4.400 727.240 1496.000 728.640 ;
        RECT 3.990 721.840 1496.000 727.240 ;
        RECT 4.400 720.440 1496.000 721.840 ;
        RECT 3.990 715.040 1496.000 720.440 ;
        RECT 4.400 713.640 1496.000 715.040 ;
        RECT 3.990 708.240 1496.000 713.640 ;
        RECT 4.400 706.840 1495.600 708.240 ;
        RECT 3.990 701.440 1496.000 706.840 ;
        RECT 4.400 700.040 1496.000 701.440 ;
        RECT 3.990 694.640 1496.000 700.040 ;
        RECT 4.400 693.240 1496.000 694.640 ;
        RECT 3.990 687.840 1496.000 693.240 ;
        RECT 4.400 686.440 1496.000 687.840 ;
        RECT 3.990 681.040 1496.000 686.440 ;
        RECT 4.400 679.640 1495.600 681.040 ;
        RECT 3.990 674.240 1496.000 679.640 ;
        RECT 4.400 672.840 1496.000 674.240 ;
        RECT 3.990 667.440 1496.000 672.840 ;
        RECT 4.400 666.040 1496.000 667.440 ;
        RECT 3.990 660.640 1496.000 666.040 ;
        RECT 4.400 659.240 1496.000 660.640 ;
        RECT 3.990 653.840 1496.000 659.240 ;
        RECT 4.400 652.440 1495.600 653.840 ;
        RECT 3.990 647.040 1496.000 652.440 ;
        RECT 4.400 645.640 1496.000 647.040 ;
        RECT 3.990 640.240 1496.000 645.640 ;
        RECT 4.400 638.840 1496.000 640.240 ;
        RECT 3.990 633.440 1496.000 638.840 ;
        RECT 4.400 632.040 1496.000 633.440 ;
        RECT 3.990 626.640 1496.000 632.040 ;
        RECT 4.400 625.240 1495.600 626.640 ;
        RECT 3.990 619.840 1496.000 625.240 ;
        RECT 4.400 618.440 1496.000 619.840 ;
        RECT 3.990 613.040 1496.000 618.440 ;
        RECT 4.400 611.640 1496.000 613.040 ;
        RECT 3.990 606.240 1496.000 611.640 ;
        RECT 4.400 604.840 1496.000 606.240 ;
        RECT 3.990 599.440 1496.000 604.840 ;
        RECT 4.400 598.040 1495.600 599.440 ;
        RECT 3.990 592.640 1496.000 598.040 ;
        RECT 4.400 591.240 1496.000 592.640 ;
        RECT 3.990 585.840 1496.000 591.240 ;
        RECT 4.400 584.440 1496.000 585.840 ;
        RECT 3.990 579.040 1496.000 584.440 ;
        RECT 4.400 577.640 1496.000 579.040 ;
        RECT 3.990 572.240 1496.000 577.640 ;
        RECT 4.400 570.840 1495.600 572.240 ;
        RECT 3.990 565.440 1496.000 570.840 ;
        RECT 4.400 564.040 1496.000 565.440 ;
        RECT 3.990 558.640 1496.000 564.040 ;
        RECT 4.400 557.240 1496.000 558.640 ;
        RECT 3.990 551.840 1496.000 557.240 ;
        RECT 4.400 550.440 1496.000 551.840 ;
        RECT 3.990 545.040 1496.000 550.440 ;
        RECT 4.400 543.640 1495.600 545.040 ;
        RECT 3.990 538.240 1496.000 543.640 ;
        RECT 4.400 536.840 1496.000 538.240 ;
        RECT 3.990 531.440 1496.000 536.840 ;
        RECT 4.400 530.040 1496.000 531.440 ;
        RECT 3.990 524.640 1496.000 530.040 ;
        RECT 4.400 523.240 1496.000 524.640 ;
        RECT 3.990 517.840 1496.000 523.240 ;
        RECT 4.400 516.440 1495.600 517.840 ;
        RECT 3.990 511.040 1496.000 516.440 ;
        RECT 4.400 509.640 1496.000 511.040 ;
        RECT 3.990 504.240 1496.000 509.640 ;
        RECT 4.400 502.840 1496.000 504.240 ;
        RECT 3.990 497.440 1496.000 502.840 ;
        RECT 4.400 496.040 1496.000 497.440 ;
        RECT 3.990 490.640 1496.000 496.040 ;
        RECT 4.400 489.240 1495.600 490.640 ;
        RECT 3.990 483.840 1496.000 489.240 ;
        RECT 4.400 482.440 1496.000 483.840 ;
        RECT 3.990 477.040 1496.000 482.440 ;
        RECT 4.400 475.640 1496.000 477.040 ;
        RECT 3.990 470.240 1496.000 475.640 ;
        RECT 4.400 468.840 1496.000 470.240 ;
        RECT 3.990 463.440 1496.000 468.840 ;
        RECT 4.400 462.040 1495.600 463.440 ;
        RECT 3.990 456.640 1496.000 462.040 ;
        RECT 4.400 455.240 1496.000 456.640 ;
        RECT 3.990 449.840 1496.000 455.240 ;
        RECT 4.400 448.440 1496.000 449.840 ;
        RECT 3.990 443.040 1496.000 448.440 ;
        RECT 4.400 441.640 1496.000 443.040 ;
        RECT 3.990 436.240 1496.000 441.640 ;
        RECT 4.400 434.840 1495.600 436.240 ;
        RECT 3.990 429.440 1496.000 434.840 ;
        RECT 4.400 428.040 1496.000 429.440 ;
        RECT 3.990 422.640 1496.000 428.040 ;
        RECT 4.400 421.240 1496.000 422.640 ;
        RECT 3.990 415.840 1496.000 421.240 ;
        RECT 4.400 414.440 1496.000 415.840 ;
        RECT 3.990 409.040 1496.000 414.440 ;
        RECT 4.400 407.640 1495.600 409.040 ;
        RECT 3.990 402.240 1496.000 407.640 ;
        RECT 4.400 400.840 1496.000 402.240 ;
        RECT 3.990 395.440 1496.000 400.840 ;
        RECT 4.400 394.040 1496.000 395.440 ;
        RECT 3.990 388.640 1496.000 394.040 ;
        RECT 4.400 387.240 1496.000 388.640 ;
        RECT 3.990 381.840 1496.000 387.240 ;
        RECT 4.400 380.440 1495.600 381.840 ;
        RECT 3.990 375.040 1496.000 380.440 ;
        RECT 4.400 373.640 1496.000 375.040 ;
        RECT 3.990 368.240 1496.000 373.640 ;
        RECT 4.400 366.840 1496.000 368.240 ;
        RECT 3.990 361.440 1496.000 366.840 ;
        RECT 4.400 360.040 1496.000 361.440 ;
        RECT 3.990 354.640 1496.000 360.040 ;
        RECT 4.400 353.240 1495.600 354.640 ;
        RECT 3.990 347.840 1496.000 353.240 ;
        RECT 4.400 346.440 1496.000 347.840 ;
        RECT 3.990 341.040 1496.000 346.440 ;
        RECT 4.400 339.640 1496.000 341.040 ;
        RECT 3.990 334.240 1496.000 339.640 ;
        RECT 4.400 332.840 1496.000 334.240 ;
        RECT 3.990 327.440 1496.000 332.840 ;
        RECT 4.400 326.040 1495.600 327.440 ;
        RECT 3.990 320.640 1496.000 326.040 ;
        RECT 4.400 319.240 1496.000 320.640 ;
        RECT 3.990 313.840 1496.000 319.240 ;
        RECT 4.400 312.440 1496.000 313.840 ;
        RECT 3.990 307.040 1496.000 312.440 ;
        RECT 4.400 305.640 1496.000 307.040 ;
        RECT 3.990 300.240 1496.000 305.640 ;
        RECT 4.400 298.840 1495.600 300.240 ;
        RECT 3.990 293.440 1496.000 298.840 ;
        RECT 4.400 292.040 1496.000 293.440 ;
        RECT 3.990 286.640 1496.000 292.040 ;
        RECT 4.400 285.240 1496.000 286.640 ;
        RECT 3.990 279.840 1496.000 285.240 ;
        RECT 4.400 278.440 1496.000 279.840 ;
        RECT 3.990 273.040 1496.000 278.440 ;
        RECT 4.400 271.640 1495.600 273.040 ;
        RECT 3.990 266.240 1496.000 271.640 ;
        RECT 4.400 264.840 1496.000 266.240 ;
        RECT 3.990 259.440 1496.000 264.840 ;
        RECT 4.400 258.040 1496.000 259.440 ;
        RECT 3.990 252.640 1496.000 258.040 ;
        RECT 4.400 251.240 1496.000 252.640 ;
        RECT 3.990 245.840 1496.000 251.240 ;
        RECT 4.400 244.440 1495.600 245.840 ;
        RECT 3.990 239.040 1496.000 244.440 ;
        RECT 4.400 237.640 1496.000 239.040 ;
        RECT 3.990 232.240 1496.000 237.640 ;
        RECT 4.400 230.840 1496.000 232.240 ;
        RECT 3.990 225.440 1496.000 230.840 ;
        RECT 4.400 224.040 1496.000 225.440 ;
        RECT 3.990 218.640 1496.000 224.040 ;
        RECT 4.400 217.240 1495.600 218.640 ;
        RECT 3.990 211.840 1496.000 217.240 ;
        RECT 4.400 210.440 1496.000 211.840 ;
        RECT 3.990 205.040 1496.000 210.440 ;
        RECT 4.400 203.640 1496.000 205.040 ;
        RECT 3.990 198.240 1496.000 203.640 ;
        RECT 4.400 196.840 1496.000 198.240 ;
        RECT 3.990 191.440 1496.000 196.840 ;
        RECT 4.400 190.040 1495.600 191.440 ;
        RECT 3.990 184.640 1496.000 190.040 ;
        RECT 4.400 183.240 1496.000 184.640 ;
        RECT 3.990 177.840 1496.000 183.240 ;
        RECT 4.400 176.440 1496.000 177.840 ;
        RECT 3.990 171.040 1496.000 176.440 ;
        RECT 4.400 169.640 1496.000 171.040 ;
        RECT 3.990 164.240 1496.000 169.640 ;
        RECT 4.400 162.840 1495.600 164.240 ;
        RECT 3.990 157.440 1496.000 162.840 ;
        RECT 4.400 156.040 1496.000 157.440 ;
        RECT 3.990 150.640 1496.000 156.040 ;
        RECT 4.400 149.240 1496.000 150.640 ;
        RECT 3.990 143.840 1496.000 149.240 ;
        RECT 4.400 142.440 1496.000 143.840 ;
        RECT 3.990 137.040 1496.000 142.440 ;
        RECT 4.400 135.640 1495.600 137.040 ;
        RECT 3.990 130.240 1496.000 135.640 ;
        RECT 4.400 128.840 1496.000 130.240 ;
        RECT 3.990 123.440 1496.000 128.840 ;
        RECT 4.400 122.040 1496.000 123.440 ;
        RECT 3.990 116.640 1496.000 122.040 ;
        RECT 4.400 115.240 1496.000 116.640 ;
        RECT 3.990 109.840 1496.000 115.240 ;
        RECT 4.400 108.440 1495.600 109.840 ;
        RECT 3.990 103.040 1496.000 108.440 ;
        RECT 4.400 101.640 1496.000 103.040 ;
        RECT 3.990 96.240 1496.000 101.640 ;
        RECT 4.400 94.840 1496.000 96.240 ;
        RECT 3.990 89.440 1496.000 94.840 ;
        RECT 4.400 88.040 1496.000 89.440 ;
        RECT 3.990 82.640 1496.000 88.040 ;
        RECT 4.400 81.240 1495.600 82.640 ;
        RECT 3.990 75.840 1496.000 81.240 ;
        RECT 4.400 74.440 1496.000 75.840 ;
        RECT 3.990 69.040 1496.000 74.440 ;
        RECT 4.400 67.640 1496.000 69.040 ;
        RECT 3.990 62.240 1496.000 67.640 ;
        RECT 4.400 60.840 1496.000 62.240 ;
        RECT 3.990 55.440 1496.000 60.840 ;
        RECT 4.400 54.040 1495.600 55.440 ;
        RECT 3.990 48.640 1496.000 54.040 ;
        RECT 4.400 47.240 1496.000 48.640 ;
        RECT 3.990 41.840 1496.000 47.240 ;
        RECT 4.400 40.440 1496.000 41.840 ;
        RECT 3.990 35.040 1496.000 40.440 ;
        RECT 4.400 33.640 1496.000 35.040 ;
        RECT 3.990 28.240 1496.000 33.640 ;
        RECT 3.990 26.840 1495.600 28.240 ;
        RECT 3.990 10.715 1496.000 26.840 ;
      LAYER met4 ;
        RECT 10.910 109.655 20.640 1176.225 ;
        RECT 23.040 109.655 97.440 1176.225 ;
        RECT 99.840 109.655 174.240 1176.225 ;
        RECT 176.640 109.655 251.040 1176.225 ;
        RECT 253.440 997.845 327.840 1176.225 ;
        RECT 330.240 997.845 404.640 1176.225 ;
        RECT 407.040 997.845 481.440 1176.225 ;
        RECT 483.840 997.845 558.240 1176.225 ;
        RECT 560.640 997.845 635.040 1176.225 ;
        RECT 637.440 997.845 711.840 1176.225 ;
        RECT 714.240 997.845 788.640 1176.225 ;
        RECT 791.040 997.845 865.440 1176.225 ;
        RECT 867.840 997.845 942.240 1176.225 ;
        RECT 253.440 310.635 942.240 997.845 ;
        RECT 253.440 109.655 327.840 310.635 ;
        RECT 330.240 109.655 404.640 310.635 ;
        RECT 407.040 109.655 481.440 310.635 ;
        RECT 483.840 109.655 558.240 310.635 ;
        RECT 560.640 109.655 635.040 310.635 ;
        RECT 637.440 109.655 711.840 310.635 ;
        RECT 714.240 109.655 788.640 310.635 ;
        RECT 791.040 109.655 865.440 310.635 ;
        RECT 867.840 109.655 942.240 310.635 ;
        RECT 944.640 109.655 1019.040 1176.225 ;
        RECT 1021.440 939.040 1095.840 1176.225 ;
        RECT 1021.440 785.440 1048.980 939.040 ;
        RECT 1051.380 922.605 1095.840 939.040 ;
        RECT 1098.240 924.680 1172.640 1176.225 ;
        RECT 1175.040 924.680 1249.440 1176.225 ;
        RECT 1098.240 922.605 1249.440 924.680 ;
        RECT 1051.380 803.195 1249.440 922.605 ;
        RECT 1051.380 785.440 1095.840 803.195 ;
        RECT 1021.440 634.400 1095.840 785.440 ;
        RECT 1021.440 486.240 1048.980 634.400 ;
        RECT 1051.380 486.240 1095.840 634.400 ;
        RECT 1021.440 362.400 1095.840 486.240 ;
        RECT 1021.440 187.040 1048.980 362.400 ;
        RECT 1051.380 347.085 1095.840 362.400 ;
        RECT 1098.240 800.440 1249.440 803.195 ;
        RECT 1098.240 619.240 1172.640 800.440 ;
        RECT 1175.040 619.240 1249.440 800.440 ;
        RECT 1098.240 499.115 1249.440 619.240 ;
        RECT 1098.240 347.085 1172.640 499.115 ;
        RECT 1175.040 347.085 1249.440 499.115 ;
        RECT 1051.380 202.515 1249.440 347.085 ;
        RECT 1051.380 187.040 1095.840 202.515 ;
        RECT 1021.440 109.655 1095.840 187.040 ;
        RECT 1098.240 109.655 1172.640 202.515 ;
        RECT 1175.040 109.655 1249.440 202.515 ;
        RECT 1251.840 109.655 1326.240 1176.225 ;
        RECT 1328.640 109.655 1403.040 1176.225 ;
        RECT 1405.440 109.655 1479.065 1176.225 ;
      LAYER met5 ;
        RECT 10.700 201.500 1244.680 1029.300 ;
  END
END aether_soc
END LIBRARY

