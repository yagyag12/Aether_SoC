// Created with Corsair v1.0.4

`ifndef __UART_REGS_VH
`define __UART_REGS_VH

`define UART_BASE_ADDR 0
`define UART_DATA_WIDTH 32
`define UART_ADDR_WIDTH 32

// UART_CTRL - UART CONTROL REGISTER
`define UART_UART_CTRL_ADDR 32'h0
`define UART_UART_CTRL_RESET 32'h0

// UART_CTRL.UART_EN - Enable Uart
`define UART_UART_CTRL_UART_EN_WIDTH 1
`define UART_UART_CTRL_UART_EN_LSB 0
`define UART_UART_CTRL_UART_EN_MASK 32'h0
`define UART_UART_CTRL_UART_EN_RESET 1'h0

// UART_CTRL.TX_EN - Enable Transmitter
`define UART_UART_CTRL_TX_EN_WIDTH 1
`define UART_UART_CTRL_TX_EN_LSB 1
`define UART_UART_CTRL_TX_EN_MASK 32'h0
`define UART_UART_CTRL_TX_EN_RESET 1'h0

// UART_CTRL.RX_EN - Enable Receiver
`define UART_UART_CTRL_RX_EN_WIDTH 1
`define UART_UART_CTRL_RX_EN_LSB 2
`define UART_UART_CTRL_RX_EN_MASK 32'h0
`define UART_UART_CTRL_RX_EN_RESET 1'h0

// UART_CTRL.TX_IRQ_EN - Enable TX Interrupt
`define UART_UART_CTRL_TX_IRQ_EN_WIDTH 1
`define UART_UART_CTRL_TX_IRQ_EN_LSB 3
`define UART_UART_CTRL_TX_IRQ_EN_MASK 32'h0
`define UART_UART_CTRL_TX_IRQ_EN_RESET 1'h0

// UART_CTRL.RX_IRQ_EN - Enable RX Interrupt
`define UART_UART_CTRL_RX_IRQ_EN_WIDTH 1
`define UART_UART_CTRL_RX_IRQ_EN_LSB 4
`define UART_UART_CTRL_RX_IRQ_EN_MASK 32'h0
`define UART_UART_CTRL_RX_IRQ_EN_RESET 1'h0

// UART_CTRL.BAUD_SEL - Baud Rate Selection (00->4800 / 01->9600 / 10->57600 / 11->115200)
`define UART_UART_CTRL_BAUD_SEL_WIDTH 2
`define UART_UART_CTRL_BAUD_SEL_LSB 5
`define UART_UART_CTRL_BAUD_SEL_MASK 32'h0
`define UART_UART_CTRL_BAUD_SEL_RESET 2'h0


// UART_STAT - UART STATUS REGISTER
`define UART_UART_STAT_ADDR 32'h4
`define UART_UART_STAT_RESET 32'h12

// UART_STAT.TX_RDY - Transmitter Ready
`define UART_UART_STAT_TX_RDY_WIDTH 1
`define UART_UART_STAT_TX_RDY_LSB 1
`define UART_UART_STAT_TX_RDY_MASK 32'h4
`define UART_UART_STAT_TX_RDY_RESET 1'h1

// UART_STAT.TX_DONE - Transmitter Done
`define UART_UART_STAT_TX_DONE_WIDTH 1
`define UART_UART_STAT_TX_DONE_LSB 2
`define UART_UART_STAT_TX_DONE_MASK 32'h4
`define UART_UART_STAT_TX_DONE_RESET 1'h0

// UART_STAT.RX_RDY - Receiver Ready
`define UART_UART_STAT_RX_RDY_WIDTH 1
`define UART_UART_STAT_RX_RDY_LSB 4
`define UART_UART_STAT_RX_RDY_MASK 32'h4
`define UART_UART_STAT_RX_RDY_RESET 1'h1

// UART_STAT.RX_DONE - Receiver Done
`define UART_UART_STAT_RX_DONE_WIDTH 1
`define UART_UART_STAT_RX_DONE_LSB 5
`define UART_UART_STAT_RX_DONE_MASK 32'h4
`define UART_UART_STAT_RX_DONE_RESET 1'h0

// UART_STAT.RX_FULL - RX Buffer Full
`define UART_UART_STAT_RX_FULL_WIDTH 1
`define UART_UART_STAT_RX_FULL_LSB 6
`define UART_UART_STAT_RX_FULL_MASK 32'h4
`define UART_UART_STAT_RX_FULL_RESET 1'h0


// UART_DATA - UART DATA REGISTER
`define UART_UART_DATA_ADDR 32'h8
`define UART_UART_DATA_RESET 32'h0

// UART_DATA.TX_DATA - UART TX Data
`define UART_UART_DATA_TX_DATA_WIDTH 8
`define UART_UART_DATA_TX_DATA_LSB 0
`define UART_UART_DATA_TX_DATA_MASK 32'h8
`define UART_UART_DATA_TX_DATA_RESET 8'h0

// UART_DATA.RX_DATA - UART RX Data
`define UART_UART_DATA_RX_DATA_WIDTH 8
`define UART_UART_DATA_RX_DATA_LSB 8
`define UART_UART_DATA_RX_DATA_MASK 32'h8
`define UART_UART_DATA_RX_DATA_RESET 8'h0


`endif // __UART_REGS_VH