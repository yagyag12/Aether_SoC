VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spi_top
  CLASS BLOCK ;
  FOREIGN spi_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.590 10.640 23.190 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 48.730 10.640 50.330 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.870 10.640 77.470 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.010 10.640 104.610 109.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 25.620 114.320 27.220 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 50.100 114.320 51.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 74.580 114.320 76.180 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 99.060 114.320 100.660 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.290 10.640 19.890 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.430 10.640 47.030 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 72.570 10.640 74.170 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.710 10.640 101.310 109.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 22.320 114.320 23.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 46.800 114.320 48.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 71.280 114.320 72.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 95.760 114.320 97.360 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END clk
  PIN i_spi_csn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END i_spi_csn
  PIN io_spi_clk
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END io_spi_clk
  PIN io_spi_miso_bit
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_spi_miso_bit
  PIN io_spi_mosi_bit
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_spi_mosi_bit
  PIN o_spi_cs[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 23.840 120.000 24.440 ;
    END
  END o_spi_cs[0]
  PIN o_spi_cs[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 20.440 120.000 21.040 ;
    END
  END o_spi_cs[1]
  PIN o_spi_cs[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 17.040 120.000 17.640 ;
    END
  END o_spi_cs[2]
  PIN o_spi_cs[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 37.440 120.000 38.040 ;
    END
  END o_spi_cs[3]
  PIN raddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 44.240 120.000 44.840 ;
    END
  END raddr[0]
  PIN raddr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 47.640 120.000 48.240 ;
    END
  END raddr[10]
  PIN raddr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 64.640 120.000 65.240 ;
    END
  END raddr[11]
  PIN raddr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 68.040 120.000 68.640 ;
    END
  END raddr[12]
  PIN raddr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 61.240 120.000 61.840 ;
    END
  END raddr[13]
  PIN raddr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 71.440 120.000 72.040 ;
    END
  END raddr[14]
  PIN raddr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 57.840 120.000 58.440 ;
    END
  END raddr[15]
  PIN raddr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 105.440 120.000 106.040 ;
    END
  END raddr[16]
  PIN raddr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 98.640 120.000 99.240 ;
    END
  END raddr[17]
  PIN raddr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 91.840 120.000 92.440 ;
    END
  END raddr[18]
  PIN raddr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 88.440 120.000 89.040 ;
    END
  END raddr[19]
  PIN raddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 34.040 120.000 34.640 ;
    END
  END raddr[1]
  PIN raddr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 108.840 120.000 109.440 ;
    END
  END raddr[20]
  PIN raddr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 112.240 120.000 112.840 ;
    END
  END raddr[21]
  PIN raddr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 115.640 120.000 116.240 ;
    END
  END raddr[22]
  PIN raddr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 102.040 120.000 102.640 ;
    END
  END raddr[23]
  PIN raddr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 85.040 120.000 85.640 ;
    END
  END raddr[24]
  PIN raddr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 30.640 120.000 31.240 ;
    END
  END raddr[25]
  PIN raddr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 119.040 120.000 119.640 ;
    END
  END raddr[26]
  PIN raddr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 95.240 120.000 95.840 ;
    END
  END raddr[27]
  PIN raddr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 78.240 120.000 78.840 ;
    END
  END raddr[28]
  PIN raddr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 0.040 120.000 0.640 ;
    END
  END raddr[29]
  PIN raddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 13.640 120.000 14.240 ;
    END
  END raddr[2]
  PIN raddr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 81.640 120.000 82.240 ;
    END
  END raddr[30]
  PIN raddr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 74.840 120.000 75.440 ;
    END
  END raddr[31]
  PIN raddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 10.240 120.000 10.840 ;
    END
  END raddr[3]
  PIN raddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 40.840 120.000 41.440 ;
    END
  END raddr[4]
  PIN raddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 6.840 120.000 7.440 ;
    END
  END raddr[5]
  PIN raddr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 54.440 120.000 55.040 ;
    END
  END raddr[6]
  PIN raddr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 51.040 120.000 51.640 ;
    END
  END raddr[7]
  PIN raddr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 3.440 120.000 4.040 ;
    END
  END raddr[8]
  PIN raddr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 116.000 27.240 120.000 27.840 ;
    END
  END raddr[9]
  PIN rdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 19.410 116.000 19.690 120.000 ;
    END
  END rdata[0]
  PIN rdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 116.000 55.110 120.000 ;
    END
  END rdata[10]
  PIN rdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 51.610 116.000 51.890 120.000 ;
    END
  END rdata[11]
  PIN rdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 116.000 74.430 120.000 ;
    END
  END rdata[12]
  PIN rdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 9.750 116.000 10.030 120.000 ;
    END
  END rdata[13]
  PIN rdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 116.000 48.670 120.000 ;
    END
  END rdata[14]
  PIN rdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 116.000 67.990 120.000 ;
    END
  END rdata[15]
  PIN rdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END rdata[16]
  PIN rdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 116.000 26.130 120.000 ;
    END
  END rdata[17]
  PIN rdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END rdata[18]
  PIN rdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END rdata[19]
  PIN rdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 116.000 61.550 120.000 ;
    END
  END rdata[1]
  PIN rdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END rdata[20]
  PIN rdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END rdata[21]
  PIN rdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END rdata[22]
  PIN rdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END rdata[23]
  PIN rdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 116.000 116.290 120.000 ;
    END
  END rdata[24]
  PIN rdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 116.000 119.510 120.000 ;
    END
  END rdata[25]
  PIN rdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END rdata[26]
  PIN rdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END rdata[27]
  PIN rdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 116.000 90.530 120.000 ;
    END
  END rdata[28]
  PIN rdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END rdata[29]
  PIN rdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.730 116.000 39.010 120.000 ;
    END
  END rdata[2]
  PIN rdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END rdata[30]
  PIN rdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END rdata[31]
  PIN rdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 116.000 71.210 120.000 ;
    END
  END rdata[3]
  PIN rdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.070 116.000 29.350 120.000 ;
    END
  END rdata[4]
  PIN rdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END rdata[5]
  PIN rdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END rdata[6]
  PIN rdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END rdata[7]
  PIN rdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 116.000 16.470 120.000 ;
    END
  END rdata[8]
  PIN rdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.170 116.000 45.450 120.000 ;
    END
  END rdata[9]
  PIN ren
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 116.000 22.910 120.000 ;
    END
  END ren
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 116.000 64.770 120.000 ;
    END
  END rst
  PIN rvalid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 6.530 116.000 6.810 120.000 ;
    END
  END rvalid
  PIN waddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END waddr[0]
  PIN waddr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 116.000 93.750 120.000 ;
    END
  END waddr[10]
  PIN waddr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3.310 116.000 3.590 120.000 ;
    END
  END waddr[11]
  PIN waddr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 116.000 80.870 120.000 ;
    END
  END waddr[12]
  PIN waddr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END waddr[13]
  PIN waddr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END waddr[14]
  PIN waddr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END waddr[15]
  PIN waddr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END waddr[16]
  PIN waddr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 116.000 100.190 120.000 ;
    END
  END waddr[17]
  PIN waddr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 116.000 84.090 120.000 ;
    END
  END waddr[18]
  PIN waddr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 116.000 87.310 120.000 ;
    END
  END waddr[19]
  PIN waddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 116.000 96.970 120.000 ;
    END
  END waddr[1]
  PIN waddr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 116.000 58.330 120.000 ;
    END
  END waddr[20]
  PIN waddr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END waddr[21]
  PIN waddr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END waddr[22]
  PIN waddr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END waddr[23]
  PIN waddr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 116.000 77.650 120.000 ;
    END
  END waddr[24]
  PIN waddr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 116.000 106.630 120.000 ;
    END
  END waddr[25]
  PIN waddr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END waddr[26]
  PIN waddr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END waddr[27]
  PIN waddr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 116.000 0.370 120.000 ;
    END
  END waddr[28]
  PIN waddr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 116.000 42.230 120.000 ;
    END
  END waddr[29]
  PIN waddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END waddr[2]
  PIN waddr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 116.000 13.250 120.000 ;
    END
  END waddr[30]
  PIN waddr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END waddr[31]
  PIN waddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END waddr[3]
  PIN waddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END waddr[4]
  PIN waddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 116.000 103.410 120.000 ;
    END
  END waddr[5]
  PIN waddr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 116.000 109.850 120.000 ;
    END
  END waddr[6]
  PIN waddr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 116.000 113.070 120.000 ;
    END
  END waddr[7]
  PIN waddr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END waddr[8]
  PIN waddr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END waddr[9]
  PIN wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wdata[0]
  PIN wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wdata[10]
  PIN wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wdata[11]
  PIN wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 116.000 35.790 120.000 ;
    END
  END wdata[12]
  PIN wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 116.000 32.570 120.000 ;
    END
  END wdata[13]
  PIN wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END wdata[14]
  PIN wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END wdata[15]
  PIN wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wdata[16]
  PIN wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wdata[17]
  PIN wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wdata[18]
  PIN wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wdata[19]
  PIN wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wdata[1]
  PIN wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wdata[20]
  PIN wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wdata[21]
  PIN wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wdata[22]
  PIN wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wdata[23]
  PIN wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wdata[24]
  PIN wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wdata[25]
  PIN wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END wdata[26]
  PIN wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wdata[27]
  PIN wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END wdata[28]
  PIN wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wdata[29]
  PIN wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END wdata[2]
  PIN wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wdata[30]
  PIN wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END wdata[31]
  PIN wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END wdata[3]
  PIN wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wdata[4]
  PIN wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wdata[5]
  PIN wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END wdata[6]
  PIN wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wdata[7]
  PIN wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wdata[8]
  PIN wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wdata[9]
  PIN wen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wen
  PIN wready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END wready
  PIN wstrb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wstrb[0]
  PIN wstrb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wstrb[1]
  PIN wstrb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END wstrb[2]
  PIN wstrb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END wstrb[3]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 114.270 108.885 ;
      LAYER li1 ;
        RECT 5.520 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 0.070 9.560 119.530 109.780 ;
      LAYER met2 ;
        RECT 0.650 115.720 3.030 119.525 ;
        RECT 3.870 115.720 6.250 119.525 ;
        RECT 7.090 115.720 9.470 119.525 ;
        RECT 10.310 115.720 12.690 119.525 ;
        RECT 13.530 115.720 15.910 119.525 ;
        RECT 16.750 115.720 19.130 119.525 ;
        RECT 19.970 115.720 22.350 119.525 ;
        RECT 23.190 115.720 25.570 119.525 ;
        RECT 26.410 115.720 28.790 119.525 ;
        RECT 29.630 115.720 32.010 119.525 ;
        RECT 32.850 115.720 35.230 119.525 ;
        RECT 36.070 115.720 38.450 119.525 ;
        RECT 39.290 115.720 41.670 119.525 ;
        RECT 42.510 115.720 44.890 119.525 ;
        RECT 45.730 115.720 48.110 119.525 ;
        RECT 48.950 115.720 51.330 119.525 ;
        RECT 52.170 115.720 54.550 119.525 ;
        RECT 55.390 115.720 57.770 119.525 ;
        RECT 58.610 115.720 60.990 119.525 ;
        RECT 61.830 115.720 64.210 119.525 ;
        RECT 65.050 115.720 67.430 119.525 ;
        RECT 68.270 115.720 70.650 119.525 ;
        RECT 71.490 115.720 73.870 119.525 ;
        RECT 74.710 115.720 77.090 119.525 ;
        RECT 77.930 115.720 80.310 119.525 ;
        RECT 81.150 115.720 83.530 119.525 ;
        RECT 84.370 115.720 86.750 119.525 ;
        RECT 87.590 115.720 89.970 119.525 ;
        RECT 90.810 115.720 93.190 119.525 ;
        RECT 94.030 115.720 96.410 119.525 ;
        RECT 97.250 115.720 99.630 119.525 ;
        RECT 100.470 115.720 102.850 119.525 ;
        RECT 103.690 115.720 106.070 119.525 ;
        RECT 106.910 115.720 109.290 119.525 ;
        RECT 110.130 115.720 112.510 119.525 ;
        RECT 113.350 115.720 115.730 119.525 ;
        RECT 116.570 115.720 118.950 119.525 ;
        RECT 0.100 4.280 119.500 115.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
      LAYER met3 ;
        RECT 4.400 118.640 115.600 119.505 ;
        RECT 3.990 116.640 116.000 118.640 ;
        RECT 4.400 115.240 115.600 116.640 ;
        RECT 3.990 113.240 116.000 115.240 ;
        RECT 4.400 111.840 115.600 113.240 ;
        RECT 3.990 109.840 116.000 111.840 ;
        RECT 4.400 108.440 115.600 109.840 ;
        RECT 3.990 106.440 116.000 108.440 ;
        RECT 4.400 105.040 115.600 106.440 ;
        RECT 3.990 103.040 116.000 105.040 ;
        RECT 4.400 101.640 115.600 103.040 ;
        RECT 3.990 99.640 116.000 101.640 ;
        RECT 4.400 98.240 115.600 99.640 ;
        RECT 3.990 96.240 116.000 98.240 ;
        RECT 4.400 94.840 115.600 96.240 ;
        RECT 3.990 92.840 116.000 94.840 ;
        RECT 4.400 91.440 115.600 92.840 ;
        RECT 3.990 89.440 116.000 91.440 ;
        RECT 4.400 88.040 115.600 89.440 ;
        RECT 3.990 86.040 116.000 88.040 ;
        RECT 4.400 84.640 115.600 86.040 ;
        RECT 3.990 82.640 116.000 84.640 ;
        RECT 4.400 81.240 115.600 82.640 ;
        RECT 3.990 79.240 116.000 81.240 ;
        RECT 4.400 77.840 115.600 79.240 ;
        RECT 3.990 75.840 116.000 77.840 ;
        RECT 4.400 74.440 115.600 75.840 ;
        RECT 3.990 72.440 116.000 74.440 ;
        RECT 4.400 71.040 115.600 72.440 ;
        RECT 3.990 69.040 116.000 71.040 ;
        RECT 4.400 67.640 115.600 69.040 ;
        RECT 3.990 65.640 116.000 67.640 ;
        RECT 4.400 64.240 115.600 65.640 ;
        RECT 3.990 62.240 116.000 64.240 ;
        RECT 4.400 60.840 115.600 62.240 ;
        RECT 3.990 58.840 116.000 60.840 ;
        RECT 4.400 57.440 115.600 58.840 ;
        RECT 3.990 55.440 116.000 57.440 ;
        RECT 4.400 54.040 115.600 55.440 ;
        RECT 3.990 52.040 116.000 54.040 ;
        RECT 4.400 50.640 115.600 52.040 ;
        RECT 3.990 48.640 116.000 50.640 ;
        RECT 4.400 47.240 115.600 48.640 ;
        RECT 3.990 45.240 116.000 47.240 ;
        RECT 4.400 43.840 115.600 45.240 ;
        RECT 3.990 41.840 116.000 43.840 ;
        RECT 4.400 40.440 115.600 41.840 ;
        RECT 3.990 38.440 116.000 40.440 ;
        RECT 4.400 37.040 115.600 38.440 ;
        RECT 3.990 35.040 116.000 37.040 ;
        RECT 4.400 33.640 115.600 35.040 ;
        RECT 3.990 31.640 116.000 33.640 ;
        RECT 4.400 30.240 115.600 31.640 ;
        RECT 3.990 28.240 116.000 30.240 ;
        RECT 4.400 26.840 115.600 28.240 ;
        RECT 3.990 24.840 116.000 26.840 ;
        RECT 4.400 23.440 115.600 24.840 ;
        RECT 3.990 21.440 116.000 23.440 ;
        RECT 4.400 20.040 115.600 21.440 ;
        RECT 3.990 18.040 116.000 20.040 ;
        RECT 4.400 16.640 115.600 18.040 ;
        RECT 3.990 14.640 116.000 16.640 ;
        RECT 4.400 13.240 115.600 14.640 ;
        RECT 3.990 11.240 116.000 13.240 ;
        RECT 4.400 9.840 115.600 11.240 ;
        RECT 3.990 7.840 116.000 9.840 ;
        RECT 4.400 6.440 115.600 7.840 ;
        RECT 3.990 4.440 116.000 6.440 ;
        RECT 3.990 3.040 115.600 4.440 ;
        RECT 3.990 1.040 116.000 3.040 ;
        RECT 3.990 0.175 115.600 1.040 ;
      LAYER met4 ;
        RECT 20.535 10.240 21.190 92.305 ;
        RECT 23.590 10.240 45.030 92.305 ;
        RECT 47.430 10.240 48.330 92.305 ;
        RECT 50.730 10.240 72.170 92.305 ;
        RECT 74.570 10.240 75.470 92.305 ;
        RECT 77.870 10.240 99.310 92.305 ;
        RECT 101.710 10.240 102.610 92.305 ;
        RECT 105.010 10.240 110.105 92.305 ;
        RECT 20.535 9.015 110.105 10.240 ;
  END
END spi_top
END LIBRARY

