// Created with Corsair v1.0.4

`ifndef __TIMER_REGS_VH
`define __TIMER_REGS_VH

`define TIMER_BASE_ADDR 0
`define TIMER_DATA_WIDTH 32
`define TIMER_ADDR_WIDTH 32

// TIMER_CTRL - TIMER CONTROL REGISTER
`define TIMER_TIMER_CTRL_ADDR 32'h0
`define TIMER_TIMER_CTRL_RESET 32'h0

// TIMER_CTRL.TMR_EN - Enable Timer
`define TIMER_TIMER_CTRL_TMR_EN_WIDTH 1
`define TIMER_TIMER_CTRL_TMR_EN_LSB 0
`define TIMER_TIMER_CTRL_TMR_EN_MASK 32'h0
`define TIMER_TIMER_CTRL_TMR_EN_RESET 1'h0

// TIMER_CTRL.PWM_EN - PWM Timer Enable
`define TIMER_TIMER_CTRL_PWM_EN_WIDTH 1
`define TIMER_TIMER_CTRL_PWM_EN_LSB 1
`define TIMER_TIMER_CTRL_PWM_EN_MASK 32'h0
`define TIMER_TIMER_CTRL_PWM_EN_RESET 1'h0

// TIMER_CTRL.TMR_DONE - Timer Done Flags
`define TIMER_TIMER_CTRL_TMR_DONE_WIDTH 1
`define TIMER_TIMER_CTRL_TMR_DONE_LSB 2
`define TIMER_TIMER_CTRL_TMR_DONE_MASK 32'h0
`define TIMER_TIMER_CTRL_TMR_DONE_RESET 1'h0


// TIMER0 - Timer0 Delay Register
`define TIMER_TIMER0_ADDR 32'h4
`define TIMER_TIMER0_RESET 32'h0

// TIMER0.DELAY - Timer Delay
`define TIMER_TIMER0_DELAY_WIDTH 32
`define TIMER_TIMER0_DELAY_LSB 0
`define TIMER_TIMER0_DELAY_MASK 32'h4
`define TIMER_TIMER0_DELAY_RESET 32'h0


// PWM0 - PWM0 Delay Register
`define TIMER_PWM0_ADDR 32'h8
`define TIMER_PWM0_RESET 32'h0

// PWM0.PERIOD - PWM0 Period
`define TIMER_PWM0_PERIOD_WIDTH 16
`define TIMER_PWM0_PERIOD_LSB 0
`define TIMER_PWM0_PERIOD_MASK 32'h8
`define TIMER_PWM0_PERIOD_RESET 16'h0

// PWM0.DUTY_CYCLE - PWM0 Duty Cycle
`define TIMER_PWM0_DUTY_CYCLE_WIDTH 16
`define TIMER_PWM0_DUTY_CYCLE_LSB 16
`define TIMER_PWM0_DUTY_CYCLE_MASK 32'h8
`define TIMER_PWM0_DUTY_CYCLE_RESET 16'h0


`endif // __TIMER_REGS_VH