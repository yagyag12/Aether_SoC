VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rv32_core
  CLASS BLOCK ;
  FOREIGN rv32_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 789.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 794.660 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 794.660 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 794.660 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 794.660 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 794.660 644.350 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 794.660 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 794.660 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 794.660 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 794.660 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 794.660 641.050 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 280.230 796.000 280.510 800.000 ;
    END
  END clk
  PIN dmem_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 705.270 796.000 705.550 800.000 ;
    END
  END dmem_addr[0]
  PIN dmem_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 698.830 796.000 699.110 800.000 ;
    END
  END dmem_addr[10]
  PIN dmem_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 682.730 796.000 683.010 800.000 ;
    END
  END dmem_addr[11]
  PIN dmem_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 679.510 796.000 679.790 800.000 ;
    END
  END dmem_addr[12]
  PIN dmem_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 673.070 796.000 673.350 800.000 ;
    END
  END dmem_addr[13]
  PIN dmem_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 524.950 796.000 525.230 800.000 ;
    END
  END dmem_addr[14]
  PIN dmem_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 534.610 796.000 534.890 800.000 ;
    END
  END dmem_addr[15]
  PIN dmem_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 650.530 796.000 650.810 800.000 ;
    END
  END dmem_addr[16]
  PIN dmem_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 631.210 796.000 631.490 800.000 ;
    END
  END dmem_addr[17]
  PIN dmem_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 528.170 796.000 528.450 800.000 ;
    END
  END dmem_addr[18]
  PIN dmem_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 676.290 796.000 676.570 800.000 ;
    END
  END dmem_addr[19]
  PIN dmem_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 653.750 796.000 654.030 800.000 ;
    END
  END dmem_addr[1]
  PIN dmem_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 695.610 796.000 695.890 800.000 ;
    END
  END dmem_addr[20]
  PIN dmem_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 286.670 796.000 286.950 800.000 ;
    END
  END dmem_addr[21]
  PIN dmem_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 289.890 796.000 290.170 800.000 ;
    END
  END dmem_addr[22]
  PIN dmem_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 312.430 796.000 312.710 800.000 ;
    END
  END dmem_addr[23]
  PIN dmem_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 293.110 796.000 293.390 800.000 ;
    END
  END dmem_addr[24]
  PIN dmem_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 489.530 796.000 489.810 800.000 ;
    END
  END dmem_addr[25]
  PIN dmem_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 309.210 796.000 309.490 800.000 ;
    END
  END dmem_addr[26]
  PIN dmem_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 322.090 796.000 322.370 800.000 ;
    END
  END dmem_addr[27]
  PIN dmem_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 479.870 796.000 480.150 800.000 ;
    END
  END dmem_addr[28]
  PIN dmem_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 457.330 796.000 457.610 800.000 ;
    END
  END dmem_addr[29]
  PIN dmem_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 495.970 796.000 496.250 800.000 ;
    END
  END dmem_addr[2]
  PIN dmem_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 399.370 796.000 399.650 800.000 ;
    END
  END dmem_addr[30]
  PIN dmem_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 466.990 796.000 467.270 800.000 ;
    END
  END dmem_addr[31]
  PIN dmem_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 521.730 796.000 522.010 800.000 ;
    END
  END dmem_addr[3]
  PIN dmem_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 473.430 796.000 473.710 800.000 ;
    END
  END dmem_addr[4]
  PIN dmem_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 505.630 796.000 505.910 800.000 ;
    END
  END dmem_addr[5]
  PIN dmem_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 689.170 796.000 689.450 800.000 ;
    END
  END dmem_addr[6]
  PIN dmem_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 499.190 796.000 499.470 800.000 ;
    END
  END dmem_addr[7]
  PIN dmem_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 702.050 796.000 702.330 800.000 ;
    END
  END dmem_addr[8]
  PIN dmem_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 685.950 796.000 686.230 800.000 ;
    END
  END dmem_addr[9]
  PIN dmem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 537.830 796.000 538.110 800.000 ;
    END
  END dmem_rdata[0]
  PIN dmem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 647.310 796.000 647.590 800.000 ;
    END
  END dmem_rdata[10]
  PIN dmem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 599.010 796.000 599.290 800.000 ;
    END
  END dmem_rdata[11]
  PIN dmem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 579.690 796.000 579.970 800.000 ;
    END
  END dmem_rdata[12]
  PIN dmem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 550.710 796.000 550.990 800.000 ;
    END
  END dmem_rdata[13]
  PIN dmem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 634.430 796.000 634.710 800.000 ;
    END
  END dmem_rdata[14]
  PIN dmem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 656.970 796.000 657.250 800.000 ;
    END
  END dmem_rdata[15]
  PIN dmem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 615.110 796.000 615.390 800.000 ;
    END
  END dmem_rdata[16]
  PIN dmem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 544.270 796.000 544.550 800.000 ;
    END
  END dmem_rdata[17]
  PIN dmem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 618.330 796.000 618.610 800.000 ;
    END
  END dmem_rdata[18]
  PIN dmem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 573.250 796.000 573.530 800.000 ;
    END
  END dmem_rdata[19]
  PIN dmem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 640.870 796.000 641.150 800.000 ;
    END
  END dmem_rdata[1]
  PIN dmem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 576.470 796.000 576.750 800.000 ;
    END
  END dmem_rdata[20]
  PIN dmem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 586.130 796.000 586.410 800.000 ;
    END
  END dmem_rdata[21]
  PIN dmem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 602.230 796.000 602.510 800.000 ;
    END
  END dmem_rdata[22]
  PIN dmem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 663.410 796.000 663.690 800.000 ;
    END
  END dmem_rdata[23]
  PIN dmem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 621.550 796.000 621.830 800.000 ;
    END
  END dmem_rdata[24]
  PIN dmem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 611.890 796.000 612.170 800.000 ;
    END
  END dmem_rdata[25]
  PIN dmem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 608.670 796.000 608.950 800.000 ;
    END
  END dmem_rdata[26]
  PIN dmem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 560.370 796.000 560.650 800.000 ;
    END
  END dmem_rdata[27]
  PIN dmem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 553.930 796.000 554.210 800.000 ;
    END
  END dmem_rdata[28]
  PIN dmem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 570.030 796.000 570.310 800.000 ;
    END
  END dmem_rdata[29]
  PIN dmem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 637.650 796.000 637.930 800.000 ;
    END
  END dmem_rdata[2]
  PIN dmem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 605.450 796.000 605.730 800.000 ;
    END
  END dmem_rdata[30]
  PIN dmem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 666.630 796.000 666.910 800.000 ;
    END
  END dmem_rdata[31]
  PIN dmem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 592.570 796.000 592.850 800.000 ;
    END
  END dmem_rdata[3]
  PIN dmem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 582.910 796.000 583.190 800.000 ;
    END
  END dmem_rdata[4]
  PIN dmem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 595.790 796.000 596.070 800.000 ;
    END
  END dmem_rdata[5]
  PIN dmem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 627.990 796.000 628.270 800.000 ;
    END
  END dmem_rdata[6]
  PIN dmem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 669.850 796.000 670.130 800.000 ;
    END
  END dmem_rdata[7]
  PIN dmem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 644.090 796.000 644.370 800.000 ;
    END
  END dmem_rdata[8]
  PIN dmem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 541.050 796.000 541.330 800.000 ;
    END
  END dmem_rdata[9]
  PIN dmem_ren
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 624.770 796.000 625.050 800.000 ;
    END
  END dmem_ren
  PIN dmem_rvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END dmem_rvalid
  PIN dmem_wdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END dmem_wdata[0]
  PIN dmem_wdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 328.530 796.000 328.810 800.000 ;
    END
  END dmem_wdata[10]
  PIN dmem_wdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 360.730 796.000 361.010 800.000 ;
    END
  END dmem_wdata[11]
  PIN dmem_wdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 338.190 796.000 338.470 800.000 ;
    END
  END dmem_wdata[12]
  PIN dmem_wdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 405.810 796.000 406.090 800.000 ;
    END
  END dmem_wdata[13]
  PIN dmem_wdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 347.850 796.000 348.130 800.000 ;
    END
  END dmem_wdata[14]
  PIN dmem_wdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 438.010 796.000 438.290 800.000 ;
    END
  END dmem_wdata[15]
  PIN dmem_wdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 354.290 796.000 354.570 800.000 ;
    END
  END dmem_wdata[16]
  PIN dmem_wdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 380.050 796.000 380.330 800.000 ;
    END
  END dmem_wdata[17]
  PIN dmem_wdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 486.310 796.000 486.590 800.000 ;
    END
  END dmem_wdata[18]
  PIN dmem_wdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END dmem_wdata[19]
  PIN dmem_wdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END dmem_wdata[1]
  PIN dmem_wdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END dmem_wdata[20]
  PIN dmem_wdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END dmem_wdata[21]
  PIN dmem_wdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END dmem_wdata[22]
  PIN dmem_wdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END dmem_wdata[23]
  PIN dmem_wdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END dmem_wdata[24]
  PIN dmem_wdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END dmem_wdata[25]
  PIN dmem_wdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 383.270 796.000 383.550 800.000 ;
    END
  END dmem_wdata[26]
  PIN dmem_wdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END dmem_wdata[27]
  PIN dmem_wdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END dmem_wdata[28]
  PIN dmem_wdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END dmem_wdata[29]
  PIN dmem_wdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END dmem_wdata[2]
  PIN dmem_wdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END dmem_wdata[30]
  PIN dmem_wdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 389.710 796.000 389.990 800.000 ;
    END
  END dmem_wdata[31]
  PIN dmem_wdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 299.550 796.000 299.830 800.000 ;
    END
  END dmem_wdata[3]
  PIN dmem_wdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END dmem_wdata[4]
  PIN dmem_wdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END dmem_wdata[5]
  PIN dmem_wdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END dmem_wdata[6]
  PIN dmem_wdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END dmem_wdata[7]
  PIN dmem_wdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 351.070 796.000 351.350 800.000 ;
    END
  END dmem_wdata[8]
  PIN dmem_wdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 367.170 796.000 367.450 800.000 ;
    END
  END dmem_wdata[9]
  PIN dmem_wen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 589.350 796.000 589.630 800.000 ;
    END
  END dmem_wen
  PIN dmem_wmask[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 563.590 796.000 563.870 800.000 ;
    END
  END dmem_wmask[0]
  PIN dmem_wmask[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 566.810 796.000 567.090 800.000 ;
    END
  END dmem_wmask[1]
  PIN dmem_wmask[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 557.150 796.000 557.430 800.000 ;
    END
  END dmem_wmask[2]
  PIN dmem_wmask[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 547.490 796.000 547.770 800.000 ;
    END
  END dmem_wmask[3]
  PIN imem_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 341.410 796.000 341.690 800.000 ;
    END
  END imem_addr[0]
  PIN imem_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 460.550 796.000 460.830 800.000 ;
    END
  END imem_addr[10]
  PIN imem_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 357.510 796.000 357.790 800.000 ;
    END
  END imem_addr[11]
  PIN imem_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 531.390 796.000 531.670 800.000 ;
    END
  END imem_addr[12]
  PIN imem_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 660.190 796.000 660.470 800.000 ;
    END
  END imem_addr[13]
  PIN imem_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 692.390 796.000 692.670 800.000 ;
    END
  END imem_addr[14]
  PIN imem_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 518.510 796.000 518.790 800.000 ;
    END
  END imem_addr[15]
  PIN imem_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 512.070 796.000 512.350 800.000 ;
    END
  END imem_addr[16]
  PIN imem_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 492.750 796.000 493.030 800.000 ;
    END
  END imem_addr[17]
  PIN imem_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 508.850 796.000 509.130 800.000 ;
    END
  END imem_addr[18]
  PIN imem_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 502.410 796.000 502.690 800.000 ;
    END
  END imem_addr[19]
  PIN imem_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 515.290 796.000 515.570 800.000 ;
    END
  END imem_addr[1]
  PIN imem_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 421.910 796.000 422.190 800.000 ;
    END
  END imem_addr[20]
  PIN imem_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 296.330 796.000 296.610 800.000 ;
    END
  END imem_addr[21]
  PIN imem_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 441.230 796.000 441.510 800.000 ;
    END
  END imem_addr[22]
  PIN imem_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 415.470 796.000 415.750 800.000 ;
    END
  END imem_addr[23]
  PIN imem_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 376.830 796.000 377.110 800.000 ;
    END
  END imem_addr[24]
  PIN imem_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 325.310 796.000 325.590 800.000 ;
    END
  END imem_addr[25]
  PIN imem_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 444.450 796.000 444.730 800.000 ;
    END
  END imem_addr[26]
  PIN imem_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 454.110 796.000 454.390 800.000 ;
    END
  END imem_addr[27]
  PIN imem_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 434.790 796.000 435.070 800.000 ;
    END
  END imem_addr[28]
  PIN imem_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 302.770 796.000 303.050 800.000 ;
    END
  END imem_addr[29]
  PIN imem_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 476.650 796.000 476.930 800.000 ;
    END
  END imem_addr[2]
  PIN imem_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 318.870 796.000 319.150 800.000 ;
    END
  END imem_addr[30]
  PIN imem_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 373.610 796.000 373.890 800.000 ;
    END
  END imem_addr[31]
  PIN imem_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 483.090 796.000 483.370 800.000 ;
    END
  END imem_addr[3]
  PIN imem_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 396.150 796.000 396.430 800.000 ;
    END
  END imem_addr[4]
  PIN imem_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 463.770 796.000 464.050 800.000 ;
    END
  END imem_addr[5]
  PIN imem_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 470.210 796.000 470.490 800.000 ;
    END
  END imem_addr[6]
  PIN imem_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 425.130 796.000 425.410 800.000 ;
    END
  END imem_addr[7]
  PIN imem_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 450.890 796.000 451.170 800.000 ;
    END
  END imem_addr[8]
  PIN imem_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 412.250 796.000 412.530 800.000 ;
    END
  END imem_addr[9]
  PIN imem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 331.750 796.000 332.030 800.000 ;
    END
  END imem_rdata[0]
  PIN imem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END imem_rdata[10]
  PIN imem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END imem_rdata[11]
  PIN imem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END imem_rdata[12]
  PIN imem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END imem_rdata[13]
  PIN imem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END imem_rdata[14]
  PIN imem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END imem_rdata[15]
  PIN imem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END imem_rdata[16]
  PIN imem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END imem_rdata[17]
  PIN imem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END imem_rdata[18]
  PIN imem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END imem_rdata[19]
  PIN imem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 344.630 796.000 344.910 800.000 ;
    END
  END imem_rdata[1]
  PIN imem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END imem_rdata[20]
  PIN imem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END imem_rdata[21]
  PIN imem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END imem_rdata[22]
  PIN imem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END imem_rdata[23]
  PIN imem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 447.670 796.000 447.950 800.000 ;
    END
  END imem_rdata[24]
  PIN imem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 796.000 428.630 800.000 ;
    END
  END imem_rdata[25]
  PIN imem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 402.590 796.000 402.870 800.000 ;
    END
  END imem_rdata[26]
  PIN imem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 431.570 796.000 431.850 800.000 ;
    END
  END imem_rdata[27]
  PIN imem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 409.030 796.000 409.310 800.000 ;
    END
  END imem_rdata[28]
  PIN imem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 315.650 796.000 315.930 800.000 ;
    END
  END imem_rdata[29]
  PIN imem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 363.950 796.000 364.230 800.000 ;
    END
  END imem_rdata[2]
  PIN imem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 386.490 796.000 386.770 800.000 ;
    END
  END imem_rdata[30]
  PIN imem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 418.690 796.000 418.970 800.000 ;
    END
  END imem_rdata[31]
  PIN imem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 370.390 796.000 370.670 800.000 ;
    END
  END imem_rdata[3]
  PIN imem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 796.000 393.210 800.000 ;
    END
  END imem_rdata[4]
  PIN imem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 334.970 796.000 335.250 800.000 ;
    END
  END imem_rdata[5]
  PIN imem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 305.990 796.000 306.270 800.000 ;
    END
  END imem_rdata[6]
  PIN imem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END imem_rdata[7]
  PIN imem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END imem_rdata[8]
  PIN imem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END imem_rdata[9]
  PIN rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 283.450 796.000 283.730 800.000 ;
    END
  END rstn
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 794.610 788.885 ;
      LAYER li1 ;
        RECT 5.520 10.795 794.420 788.885 ;
      LAYER met1 ;
        RECT 4.210 10.640 794.420 789.040 ;
      LAYER met2 ;
        RECT 4.230 795.720 279.950 796.690 ;
        RECT 280.790 795.720 283.170 796.690 ;
        RECT 284.010 795.720 286.390 796.690 ;
        RECT 287.230 795.720 289.610 796.690 ;
        RECT 290.450 795.720 292.830 796.690 ;
        RECT 293.670 795.720 296.050 796.690 ;
        RECT 296.890 795.720 299.270 796.690 ;
        RECT 300.110 795.720 302.490 796.690 ;
        RECT 303.330 795.720 305.710 796.690 ;
        RECT 306.550 795.720 308.930 796.690 ;
        RECT 309.770 795.720 312.150 796.690 ;
        RECT 312.990 795.720 315.370 796.690 ;
        RECT 316.210 795.720 318.590 796.690 ;
        RECT 319.430 795.720 321.810 796.690 ;
        RECT 322.650 795.720 325.030 796.690 ;
        RECT 325.870 795.720 328.250 796.690 ;
        RECT 329.090 795.720 331.470 796.690 ;
        RECT 332.310 795.720 334.690 796.690 ;
        RECT 335.530 795.720 337.910 796.690 ;
        RECT 338.750 795.720 341.130 796.690 ;
        RECT 341.970 795.720 344.350 796.690 ;
        RECT 345.190 795.720 347.570 796.690 ;
        RECT 348.410 795.720 350.790 796.690 ;
        RECT 351.630 795.720 354.010 796.690 ;
        RECT 354.850 795.720 357.230 796.690 ;
        RECT 358.070 795.720 360.450 796.690 ;
        RECT 361.290 795.720 363.670 796.690 ;
        RECT 364.510 795.720 366.890 796.690 ;
        RECT 367.730 795.720 370.110 796.690 ;
        RECT 370.950 795.720 373.330 796.690 ;
        RECT 374.170 795.720 376.550 796.690 ;
        RECT 377.390 795.720 379.770 796.690 ;
        RECT 380.610 795.720 382.990 796.690 ;
        RECT 383.830 795.720 386.210 796.690 ;
        RECT 387.050 795.720 389.430 796.690 ;
        RECT 390.270 795.720 392.650 796.690 ;
        RECT 393.490 795.720 395.870 796.690 ;
        RECT 396.710 795.720 399.090 796.690 ;
        RECT 399.930 795.720 402.310 796.690 ;
        RECT 403.150 795.720 405.530 796.690 ;
        RECT 406.370 795.720 408.750 796.690 ;
        RECT 409.590 795.720 411.970 796.690 ;
        RECT 412.810 795.720 415.190 796.690 ;
        RECT 416.030 795.720 418.410 796.690 ;
        RECT 419.250 795.720 421.630 796.690 ;
        RECT 422.470 795.720 424.850 796.690 ;
        RECT 425.690 795.720 428.070 796.690 ;
        RECT 428.910 795.720 431.290 796.690 ;
        RECT 432.130 795.720 434.510 796.690 ;
        RECT 435.350 795.720 437.730 796.690 ;
        RECT 438.570 795.720 440.950 796.690 ;
        RECT 441.790 795.720 444.170 796.690 ;
        RECT 445.010 795.720 447.390 796.690 ;
        RECT 448.230 795.720 450.610 796.690 ;
        RECT 451.450 795.720 453.830 796.690 ;
        RECT 454.670 795.720 457.050 796.690 ;
        RECT 457.890 795.720 460.270 796.690 ;
        RECT 461.110 795.720 463.490 796.690 ;
        RECT 464.330 795.720 466.710 796.690 ;
        RECT 467.550 795.720 469.930 796.690 ;
        RECT 470.770 795.720 473.150 796.690 ;
        RECT 473.990 795.720 476.370 796.690 ;
        RECT 477.210 795.720 479.590 796.690 ;
        RECT 480.430 795.720 482.810 796.690 ;
        RECT 483.650 795.720 486.030 796.690 ;
        RECT 486.870 795.720 489.250 796.690 ;
        RECT 490.090 795.720 492.470 796.690 ;
        RECT 493.310 795.720 495.690 796.690 ;
        RECT 496.530 795.720 498.910 796.690 ;
        RECT 499.750 795.720 502.130 796.690 ;
        RECT 502.970 795.720 505.350 796.690 ;
        RECT 506.190 795.720 508.570 796.690 ;
        RECT 509.410 795.720 511.790 796.690 ;
        RECT 512.630 795.720 515.010 796.690 ;
        RECT 515.850 795.720 518.230 796.690 ;
        RECT 519.070 795.720 521.450 796.690 ;
        RECT 522.290 795.720 524.670 796.690 ;
        RECT 525.510 795.720 527.890 796.690 ;
        RECT 528.730 795.720 531.110 796.690 ;
        RECT 531.950 795.720 534.330 796.690 ;
        RECT 535.170 795.720 537.550 796.690 ;
        RECT 538.390 795.720 540.770 796.690 ;
        RECT 541.610 795.720 543.990 796.690 ;
        RECT 544.830 795.720 547.210 796.690 ;
        RECT 548.050 795.720 550.430 796.690 ;
        RECT 551.270 795.720 553.650 796.690 ;
        RECT 554.490 795.720 556.870 796.690 ;
        RECT 557.710 795.720 560.090 796.690 ;
        RECT 560.930 795.720 563.310 796.690 ;
        RECT 564.150 795.720 566.530 796.690 ;
        RECT 567.370 795.720 569.750 796.690 ;
        RECT 570.590 795.720 572.970 796.690 ;
        RECT 573.810 795.720 576.190 796.690 ;
        RECT 577.030 795.720 579.410 796.690 ;
        RECT 580.250 795.720 582.630 796.690 ;
        RECT 583.470 795.720 585.850 796.690 ;
        RECT 586.690 795.720 589.070 796.690 ;
        RECT 589.910 795.720 592.290 796.690 ;
        RECT 593.130 795.720 595.510 796.690 ;
        RECT 596.350 795.720 598.730 796.690 ;
        RECT 599.570 795.720 601.950 796.690 ;
        RECT 602.790 795.720 605.170 796.690 ;
        RECT 606.010 795.720 608.390 796.690 ;
        RECT 609.230 795.720 611.610 796.690 ;
        RECT 612.450 795.720 614.830 796.690 ;
        RECT 615.670 795.720 618.050 796.690 ;
        RECT 618.890 795.720 621.270 796.690 ;
        RECT 622.110 795.720 624.490 796.690 ;
        RECT 625.330 795.720 627.710 796.690 ;
        RECT 628.550 795.720 630.930 796.690 ;
        RECT 631.770 795.720 634.150 796.690 ;
        RECT 634.990 795.720 637.370 796.690 ;
        RECT 638.210 795.720 640.590 796.690 ;
        RECT 641.430 795.720 643.810 796.690 ;
        RECT 644.650 795.720 647.030 796.690 ;
        RECT 647.870 795.720 650.250 796.690 ;
        RECT 651.090 795.720 653.470 796.690 ;
        RECT 654.310 795.720 656.690 796.690 ;
        RECT 657.530 795.720 659.910 796.690 ;
        RECT 660.750 795.720 663.130 796.690 ;
        RECT 663.970 795.720 666.350 796.690 ;
        RECT 667.190 795.720 669.570 796.690 ;
        RECT 670.410 795.720 672.790 796.690 ;
        RECT 673.630 795.720 676.010 796.690 ;
        RECT 676.850 795.720 679.230 796.690 ;
        RECT 680.070 795.720 682.450 796.690 ;
        RECT 683.290 795.720 685.670 796.690 ;
        RECT 686.510 795.720 688.890 796.690 ;
        RECT 689.730 795.720 692.110 796.690 ;
        RECT 692.950 795.720 695.330 796.690 ;
        RECT 696.170 795.720 698.550 796.690 ;
        RECT 699.390 795.720 701.770 796.690 ;
        RECT 702.610 795.720 704.990 796.690 ;
        RECT 705.830 795.720 793.910 796.690 ;
        RECT 4.230 4.280 793.910 795.720 ;
        RECT 4.230 4.000 305.710 4.280 ;
        RECT 306.550 4.000 341.130 4.280 ;
        RECT 341.970 4.000 354.010 4.280 ;
        RECT 354.850 4.000 793.910 4.280 ;
      LAYER met3 ;
        RECT 3.990 531.440 793.930 788.965 ;
        RECT 4.400 530.040 793.930 531.440 ;
        RECT 3.990 528.040 793.930 530.040 ;
        RECT 4.400 526.640 793.930 528.040 ;
        RECT 3.990 524.640 793.930 526.640 ;
        RECT 4.400 523.240 793.930 524.640 ;
        RECT 3.990 521.240 793.930 523.240 ;
        RECT 4.400 519.840 793.930 521.240 ;
        RECT 3.990 517.840 793.930 519.840 ;
        RECT 4.400 516.440 793.930 517.840 ;
        RECT 3.990 514.440 793.930 516.440 ;
        RECT 4.400 513.040 793.930 514.440 ;
        RECT 3.990 511.040 793.930 513.040 ;
        RECT 4.400 509.640 793.930 511.040 ;
        RECT 3.990 507.640 793.930 509.640 ;
        RECT 4.400 506.240 793.930 507.640 ;
        RECT 3.990 504.240 793.930 506.240 ;
        RECT 4.400 502.840 793.930 504.240 ;
        RECT 3.990 500.840 793.930 502.840 ;
        RECT 4.400 499.440 793.930 500.840 ;
        RECT 3.990 497.440 793.930 499.440 ;
        RECT 4.400 496.040 793.930 497.440 ;
        RECT 3.990 494.040 793.930 496.040 ;
        RECT 4.400 492.640 793.930 494.040 ;
        RECT 3.990 490.640 793.930 492.640 ;
        RECT 4.400 489.240 793.930 490.640 ;
        RECT 3.990 487.240 793.930 489.240 ;
        RECT 4.400 485.840 793.930 487.240 ;
        RECT 3.990 483.840 793.930 485.840 ;
        RECT 4.400 482.440 793.930 483.840 ;
        RECT 3.990 480.440 793.930 482.440 ;
        RECT 4.400 479.040 793.930 480.440 ;
        RECT 3.990 477.040 793.930 479.040 ;
        RECT 4.400 475.640 793.930 477.040 ;
        RECT 3.990 473.640 793.930 475.640 ;
        RECT 4.400 472.240 793.930 473.640 ;
        RECT 3.990 470.240 793.930 472.240 ;
        RECT 4.400 468.840 793.930 470.240 ;
        RECT 3.990 466.840 793.930 468.840 ;
        RECT 4.400 465.440 793.930 466.840 ;
        RECT 3.990 463.440 793.930 465.440 ;
        RECT 4.400 462.040 793.930 463.440 ;
        RECT 3.990 460.040 793.930 462.040 ;
        RECT 4.400 458.640 793.930 460.040 ;
        RECT 3.990 456.640 793.930 458.640 ;
        RECT 4.400 455.240 793.930 456.640 ;
        RECT 3.990 453.240 793.930 455.240 ;
        RECT 4.400 451.840 793.930 453.240 ;
        RECT 3.990 449.840 793.930 451.840 ;
        RECT 4.400 448.440 793.930 449.840 ;
        RECT 3.990 446.440 793.930 448.440 ;
        RECT 4.400 445.040 793.930 446.440 ;
        RECT 3.990 443.040 793.930 445.040 ;
        RECT 4.400 441.640 793.930 443.040 ;
        RECT 3.990 439.640 793.930 441.640 ;
        RECT 4.400 438.240 793.930 439.640 ;
        RECT 3.990 436.240 793.930 438.240 ;
        RECT 4.400 434.840 793.930 436.240 ;
        RECT 3.990 432.840 793.930 434.840 ;
        RECT 4.400 431.440 793.930 432.840 ;
        RECT 3.990 429.440 793.930 431.440 ;
        RECT 4.400 428.040 793.930 429.440 ;
        RECT 3.990 426.040 793.930 428.040 ;
        RECT 4.400 424.640 793.930 426.040 ;
        RECT 3.990 10.715 793.930 424.640 ;
      LAYER met4 ;
        RECT 133.270 120.535 174.240 787.945 ;
        RECT 176.640 120.535 177.540 787.945 ;
        RECT 179.940 120.535 327.840 787.945 ;
        RECT 330.240 120.535 331.140 787.945 ;
        RECT 333.540 120.535 481.440 787.945 ;
        RECT 483.840 120.535 484.740 787.945 ;
        RECT 487.140 120.535 635.040 787.945 ;
        RECT 637.440 120.535 638.340 787.945 ;
        RECT 640.740 120.535 656.090 787.945 ;
      LAYER met5 ;
        RECT 133.060 492.770 656.300 634.900 ;
        RECT 133.060 339.590 656.300 484.670 ;
        RECT 133.060 186.410 656.300 331.490 ;
        RECT 133.060 130.100 656.300 178.310 ;
  END
END rv32_core
END LIBRARY

