// Created with Corsair v1.0.4

`ifndef __SPI_REGS_VH
`define __SPI_REGS_VH

`define SPI_BASE_ADDR 0
`define SPI_DATA_WIDTH 32
`define SPI_ADDR_WIDTH 32

// SPI_CTRL - SPI CONTROL REGISTER
`define SPI_SPI_CTRL_ADDR 32'h0
`define SPI_SPI_CTRL_RESET 32'h0

// SPI_CTRL.SPI_EN - Enable SPI
`define SPI_SPI_CTRL_SPI_EN_WIDTH 1
`define SPI_SPI_CTRL_SPI_EN_LSB 0
`define SPI_SPI_CTRL_SPI_EN_MASK 32'h0
`define SPI_SPI_CTRL_SPI_EN_RESET 1'h0

// SPI_CTRL.MASTER_EN - Enable SPI as Master (0 -> Slave / 1 -> Master)
`define SPI_SPI_CTRL_MASTER_EN_WIDTH 1
`define SPI_SPI_CTRL_MASTER_EN_LSB 1
`define SPI_SPI_CTRL_MASTER_EN_MASK 32'h0
`define SPI_SPI_CTRL_MASTER_EN_RESET 1'h0

// SPI_CTRL.CPOL - Clock Polarity
`define SPI_SPI_CTRL_CPOL_WIDTH 1
`define SPI_SPI_CTRL_CPOL_LSB 2
`define SPI_SPI_CTRL_CPOL_MASK 32'h0
`define SPI_SPI_CTRL_CPOL_RESET 1'h0

// SPI_CTRL.CPHA - Clock Phase
`define SPI_SPI_CTRL_CPHA_WIDTH 1
`define SPI_SPI_CTRL_CPHA_LSB 3
`define SPI_SPI_CTRL_CPHA_MASK 32'h0
`define SPI_SPI_CTRL_CPHA_RESET 1'h0

// SPI_CTRL.CLK_DIV - Clock Divider for SPI Clock Generation
`define SPI_SPI_CTRL_CLK_DIV_WIDTH 8
`define SPI_SPI_CTRL_CLK_DIV_LSB 4
`define SPI_SPI_CTRL_CLK_DIV_MASK 32'h0
`define SPI_SPI_CTRL_CLK_DIV_RESET 8'h0

// SPI_CTRL.CS - Chip Select
`define SPI_SPI_CTRL_CS_WIDTH 2
`define SPI_SPI_CTRL_CS_LSB 12
`define SPI_SPI_CTRL_CS_MASK 32'h0
`define SPI_SPI_CTRL_CS_RESET 2'h0


// SPI_STAT - SPI STATUS REGISTER
`define SPI_SPI_STAT_ADDR 32'h4
`define SPI_SPI_STAT_RESET 32'h5

// SPI_STAT.TX_RDY - Transmitter Ready
`define SPI_SPI_STAT_TX_RDY_WIDTH 1
`define SPI_SPI_STAT_TX_RDY_LSB 0
`define SPI_SPI_STAT_TX_RDY_MASK 32'h4
`define SPI_SPI_STAT_TX_RDY_RESET 1'h1

// SPI_STAT.TX_DONE - Transmitter Done
`define SPI_SPI_STAT_TX_DONE_WIDTH 1
`define SPI_SPI_STAT_TX_DONE_LSB 1
`define SPI_SPI_STAT_TX_DONE_MASK 32'h4
`define SPI_SPI_STAT_TX_DONE_RESET 1'h0

// SPI_STAT.RX_RDY - Receiver Ready
`define SPI_SPI_STAT_RX_RDY_WIDTH 1
`define SPI_SPI_STAT_RX_RDY_LSB 2
`define SPI_SPI_STAT_RX_RDY_MASK 32'h4
`define SPI_SPI_STAT_RX_RDY_RESET 1'h1

// SPI_STAT.RX_DONE - Receiver Done
`define SPI_SPI_STAT_RX_DONE_WIDTH 1
`define SPI_SPI_STAT_RX_DONE_LSB 3
`define SPI_SPI_STAT_RX_DONE_MASK 32'h4
`define SPI_SPI_STAT_RX_DONE_RESET 1'h0

// SPI_STAT.BUSY - SPI is busy
`define SPI_SPI_STAT_BUSY_WIDTH 1
`define SPI_SPI_STAT_BUSY_LSB 4
`define SPI_SPI_STAT_BUSY_MASK 32'h4
`define SPI_SPI_STAT_BUSY_RESET 1'h0


// SPI_DATA - SPI DATA REGISTER
`define SPI_SPI_DATA_ADDR 32'h8
`define SPI_SPI_DATA_RESET 32'h0

// SPI_DATA.TX_DATA - SPI TX Data
`define SPI_SPI_DATA_TX_DATA_WIDTH 8
`define SPI_SPI_DATA_TX_DATA_LSB 0
`define SPI_SPI_DATA_TX_DATA_MASK 32'h8
`define SPI_SPI_DATA_TX_DATA_RESET 8'h0

// SPI_DATA.RX_DATA - SPI RX Data
`define SPI_SPI_DATA_RX_DATA_WIDTH 8
`define SPI_SPI_DATA_RX_DATA_LSB 8
`define SPI_SPI_DATA_RX_DATA_MASK 32'h8
`define SPI_SPI_DATA_RX_DATA_RESET 8'h0


`endif // __SPI_REGS_VH